//Test Bench for Floating Point Adder

`timescale 1ns/1ps

module FLOATING_POINT_ADDER_TEST_BENCH;
	reg[31:0] in1, in2;
	wire[31:0] out;

	FLOATING_POINT_ADDER_DATA_PATH DUT(in1, in2, out);

	initial begin
		$dumpfile("FLOATING_POINT_ADDER_DATA_PATH.vcd");
		$dumpvars(0, FLOATING_POINT_ADDER_TEST_BENCH);
		$monitor("%32b", DUT.out);
		//in1 = 32'b00111111100110011001100110011001;
		//in2 = 32'b00111110010011001100110011001100;
		//in1 = 32'b10111111100110011001100110011001;
		//in2 = 32'b00111110110011001100110011001100;
		in1 = 32'b10111111010011001100110011001101;                //in1 = -0.8
		in2 = 32'b10111111000110011001100110011010;		   //in2 = 0.6
	end
endmodule
